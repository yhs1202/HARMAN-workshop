package hm_pkg;
import uvm_pkg::*;
`include "3_my_seq_item.sv"
`include "4_sequence.sv"
`include "5_sequencer.sv"
`include "6_driver.sv"
`include "7_monitor.sv"
`include "8_scoreboard.sv"
`include "9_agent.sv"
`include "10_env.sv"
`include "11_test.sv"
`include "uvm_macros.svh"
    
endpackage