
interface dut_if;
    logic clock, en;
    logic [3:0] a, b;
    logic [4:0] sum;
endinterface
