`include "top.v"
`include "single_port_ram.v"
`include "line_buf_ctrl.v"
